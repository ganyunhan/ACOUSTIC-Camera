//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.08
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Sat Oct 22 12:49:41 2022

module ram5_512 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [8:0] ada;
input [15:0] din;
input [8:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[8:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({gw_gnd,adb[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h01B801C401980187011A00B60050006BFFCCFF7AFF04FF44FF0AFFA6FF46FFFB;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFE25FDEEFD14FCC4FD27FE0CFF45011C023D02CB02990296023C022F0225021C;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFDD0FDD8FDC4FD97FD98FDD0FE51FF1FFF99FFE1FF9AFF62FECEFE44FE43FE38;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h01C701A5018F020C028102AD02B70258021501CA00FC003EFF10FE5AFE13FDE0;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h03E3038A023900CBFF2CFDA2FCD0FD34FE66FFE0010F0158018301E001F80206;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hF8AFF6ABF524F4A0F53FF6D6F8F6FC0AFF23013F0286033203A503B503CB03DD;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h01A60455068E07BA090A09E50A720A90096D088E06D103CA0161FF1EFCFBFB06;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFDFBFF2A009701D202680242010EFF0EFD21FB2EF950F89BF89AF98EFBF9FED8;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFD35FE1BFF1FFF82006B015D018501B801910098FFD4FEB3FD68FCACFC94FD04;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h08BD07540630049502E40110FFB2FE6BFD37FC7FFB8FFAC9FB0FFBC2FC2AFC8C;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFED2FEA8FE22FD51FC79FC97FD50FE82001A022903CF0668085409BA0A3109ED;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h03C5044D047E048202DF000DFDACFBE1FA40F925F8A5F87BF907FA7FFBE0FDC2;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h0189017C020E02CF033D0395036D033402F3020501260093004F00B701BB02AB;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hF99DFA27FACFFBCAFDECFF7E004300AF00E40125015201D10208019C01730172;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFFBB0053FFA0FF62FF8FFF40FF1DFF0AFE8FFE2EFE0EFEA6FF57FEF2FDAFFB49;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h06C707860802085A072B051E0202FE93FB5AF8C1F82DF885F963FAD2FCA8FE39;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hF84DF76AF789F849FA6CFD3F000002560422055E07A4094209A4094B086806EA;
defparam sdpb_inst_0.INIT_RAM_11 = 256'hF961F8C9F973FB46FD48FFB501C6032704520492034000FFFEA5FCE4FAEDF9A8;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h0BD60D110D6F0C070A220784060D04F7027700F5FF58FDEAFD1FFC13FA5EF95B;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h00B202130316030A00F2FE00FAB6F744F4ABF44BF5BAF94EFE7C02F307430A7B;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFF54FE93FDFFFDD2FE19FD8AFCB7FC09FB25FABEFBCBFC78FC82FD68FE40FF40;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h08B9053C025FFFAEFD19FAF9FA81FB5CFC80FDFCFF1FFF33FED5FECBFF69FFAD;
defparam sdpb_inst_0.INIT_RAM_16 = 256'hFDBEFC02FA36FA2CFB29FD4BFF7D0175038506ED0A550D860F2F0EC00CD10ADD;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h00A90161011D011E00D5FF78FCC0F9DBF805F7DFFA11FD8B009C02560174FFB3;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h0E940E4A0DDB0C7209AB065D029FFF49FC29F931F6F5F637F778FAA8FD59FF3B;
defparam sdpb_inst_0.INIT_RAM_19 = 256'hF95DF74AF3FFF0ECEEA4EFC3F37AF818FDEF02B3074509770AE10B3B0BAA0D52;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hFEF8FFEFFFB6FFEE004B00D9027703AC048D05DA05BA045901EFFE86FC3FFAEF;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h0B030A1508BA06200294FD98F82FF374F0D4EFF9F15AF3C4F655FA04FC80FDB4;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hF8FFFD1E010202AC041506CD0A290DC70FFB0EA00C2E0A670A410B530BFC0B6F;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h029C001EFCBAFA34F969F9BDFACDFB61FBCEFB3CFA20F890F744F565F483F5B4;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h0E080B7E07E9036A00DDFF7FFF57FFC2012201EB0148FECBFC7CFC6CFE620169;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h00000000FC52F85DF8AEF717F7D6F7C8FA1DFDF002DF07690BAF0E2410190FDE;

endmodule //ram5_512
