//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Sat Oct 08 22:11:46 2022

module ram1_512 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [8:0] ada;
input [15:0] din;
input [8:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[8:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({gw_gnd,adb[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFFF1FFF7FFBBFFB1FFE1FFEA000A0041001A000A002DFFFDFFD70003FFE90005;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFFDDFFB9FFCEFFBAFFDB0010FFF5000A0013FFCAFFCC000BFFFB0004000EFFEF;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFFF90002FFD10039FFABFF66FFEFFFD7FFC4FFEAFFE100030037002E000C001B;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hFFD9002500000008FFFFFFB0FFE4FFF8002A0037002700430023FFE1FFF0FFE3;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hFFCAFFDF0002FFDAFFCEFFF1001000010001FFF6FFCCFFD8FFFBFFE6000C0002;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h000D00070019002E000DFFF40002FFCAFFD10027000CFFEB000DFFD2FFBEFFE1;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hFFFFFFD4FFEAFFD8FFC4FFD7FFF9001B000F00030006FFEEFFEBFFEAFFE3FFFA;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFFE10016FFF900160028FFF800390036FFD7FFE0FFE1FFD5002400590058003E;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h0043000BFFFEFFC4FFB0FFE3FFD6FFF0003B002C004F0055FFEDFFCCFFD5FFA8;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h001C0009FFE2FFFBFFFF001300260000FFE2FFE9FFC2FFBEFFF2FFF2FFF40038;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h000B0002000D00320007FFE4FFE1FFDAFFE0FFEDFFE0FFE6FFE7FFEDFFDFFFF0;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hFFE3000EFFC9FFBA001000120006002BFFF2FFE00001FFC7FFCB0017FFECFFD8;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFFE2FFD4FFF5FFF1FFDF00120002FFBFFFDCFFDDFFEB003000150007001DFFE2;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hFFF3001D000E0012FFE4FFD3FFF4FFF6FFE8FFFDFFF6FFF200080000FFEFFFEF;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h0004FFE300060007FFEF000AFFE7FFF5001CFFF3FFF00008FFD6FFE8FFE4FFB9;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hFFD0FFF2FFF8FFFF0027FFF0FFC80004FFF9FFEA00130008000E0014FFD7FFF8;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hFFF1FFCFFFE500160008000E0033000BFFFE0020FFEDFFF6FFE8FF9CFFCEFFF5;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h000A002CFFFFFFD3FFE1FFE7FFFA00270021000D0015FFEFFFDDFFFCFFE4FFDE;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFF5001DFFF6FFF3000EFFECFFE2FFFF000F00110010000DFFFDFFF1FFDFFFDA;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hFFED0016001FFFF3FFE4FFF8000E001B0008FFE7FFCFFFE3FFDFFFEBFFFEFFE6;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFFFEFFEAFFFB003B0004FFE50002FFBAFFCEFFFDFFE200050027001100210007;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hFFEEFFD4FFE5FFE100020016000700090007FFE6001B0014FFE900240016FFD6;
defparam sdpb_inst_0.INIT_RAM_16 = 256'hFFE1FFFDFFF90008001EFFF0FFDAFFDCFFDA0009003A001800070008000E0010;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hFFFCFFF00005FFD4FFDA0033002E000A001E000D000B002F000AFFF60011FFF4;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h001100090007001C002600140014FFF8FFDD000C000DFFF10026FFFDFFC5FFFE;
defparam sdpb_inst_0.INIT_RAM_19 = 256'hFFD1FFDFFFE5FFEC000FFFF0FFE60001FFF7FFF90018FFFFFFFFFFFBFFDFFFEF;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h00090010FFE4FFD0FFEDFFEE0003001F0019000E0019000D0021001F0006FFE0;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h001EFFFCFFE2FFDBFFD9001100390012000BFFFCFFD8FFD9FFD7FFE5000AFFFE;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hFFE4FFC8FFC6000C000DFFDDFFEDFFF9FFF2000E0008FFE9FFFC000EFFFD000E;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFFFDFFF8000B00120014000AFFE5FFD5FFD8FFE200050008FFF4000B00270002;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h000900110019FFF7FFEDFFD9FFC3FFD5FFD6FFC9FFFC0011000BFFFBFFD3FFDB;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hFFFE0020FFE9FFEAFFFFFFD6FFE500040009002E0026FFF5FFFDFFFEFFF8000C;

endmodule //ram1_512
