//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Sun Oct 09 16:33:50 2022

module ram1_512 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [8:0] ada;
input [15:0] din;
input [8:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[8:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({gw_gnd,adb[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFFD1FFBE00490015FFF1FFE5FFAA002D006FFFEEFFAFFFAD0066011E0014FFA6;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h00A4001DFF81000CFF91FF95007A0024001D00FA005C001700DA005BFFE20040;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFE1501F70143FA5902400189FF2301B7FC1FFFC40330FEF7FEFBFF9E00E30110;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hFF8801BCFE37FE5902C1018BFEBCFEDA01D500650035015DFF3900300022FFDE;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h008DFFDAFF7F0218FF6CFEF9FFE1FE3500C2FF34FCDB019D0282FF030006008F;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hFFC80052004EFEC9FF9D01550043FF1D002C001B0103014FFE3DFE7D00D0FFDB;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h001B00B3007C0018FF28FFCB00B4FFE2FFFEFFBEFEDAFF7EFFC4FEB4FF2A0068;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFF0C0067FFAEFED0FFFAFF6CFFFAFF26FED6008D007E005F0061FFE6FF6EFF43;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFFCAFFEB00230003FF93005CFF96FFAB00A2FFEE001AFFA2FFC0FF77FF61FFEE;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFFBEFF680010FFC7FF72000D0021FF23FFE70070FF31FFAC001FFFB2FFE5FF95;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFFBBFFA3FFD4004F0026FF67FF7BFFDDFFE0001A0031FF930056007BFF770010;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hFFFC000AFFB2FF9EFFE4005D000FFF7BFFB900A301290019FF3B002000F5006B;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFF64FFA90031FFD3FFCEFFDB00060060007200CA0088FFFAFFACFFE90031FFC9;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h0029001B001E0049001400120009001F003EFFC40029008900360037000DFFB8;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFF8400580069FFE1FF84FFB100870045FF860000006000A7004AFF950009004D;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hFFD4000EFFD8FF6DFF3E001300A200DB0093FFA5FFCB006700E400F8FFAAFEE1;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hFE93FF550080005CFFDAFFEA00BB013700B3FFE5002900C6004FFFD1FF9DFF5D;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h009A0020FF8BFFE3001E003C007B00BD01450116000FFF9FFFFF00660075FF9D;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFF8FFEE0011FFF0FFD0FF9BFFF70060000DFFB3008C015C008BFF78FF52FFF2;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h00380048FFA2FF4BFF8CFFE7000CFFB2FFAF0042008A0090002BFFE6008100A5;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFFF9000CFFF6FF84FEF1FEDEFF34FFCE007AFFEDFFC700AD00E200A30014FFC6;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h006C00AE0015FF7BFF33FF66FFCEFF84FF5BFFADFFC200800141010100D8006A;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h00310068008EFFC0FEECFFFB00EC00C70038FEEFFF6500D600B8002EFFACFF93;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h009CFFCEFF81000800D30077FFDDFFE4FFB9FFBFFFD4FFD80054003EFFA1FFC0;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hFF6A00370097004DFF79FED4FFDC010200900002FFC1FFD5003BFFBCFF7F0083;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h00680004FEF1FF5D00960072FFC1FF13FF6900C9008AFF7FFFBA0056003AFF7D;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h003A005FFFD6FF62FFFF00420026000BFF83FFAE00250015FFFB0004003B004A;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hFF6FFF8F002000930042FFCDFFE0FFD1FFBAFFDE001C005BFFD8FF50FFBF0026;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h00110026FFFBFF68FFB1004FFFF9FFFD0041004E0034FF81FF93004C003FFFC9;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFFDCFFBCFF8DFFBBFFDD004B0064FFF30017006BFFF6FFC3002E0015FF99FFC3;
defparam sdpb_inst_0.INIT_RAM_1E = 256'hFFBCFFC9000A0018005CFFCFFFC8009C0021FFEE0033FF74FFBF0037FF37FF1B;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hFFA6006200DF0097002000180000FFA9FF79FFD40015FF7BFF22FF57FFD00012;

endmodule //ram1_512
