//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Tue Sep 27 23:12:36 2022

module ram1_512 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [8:0] ada;
input [15:0] din;
input [8:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[8:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({gw_gnd,adb[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h0192015C00F000770065002CFFA3FF37FF21FF21FF52FF7FFF91FFB5FFD3FFE5;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFCD8FCD8FD8CFE7F001F01B6029702BB02970273022B022B022B01EC01B601B6;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFDB0FD8CFDB0FDF8FEB5FF5BFFCAFFCAFF7FFF2EFE7FFE37FE49FE25FE25FD8C;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h01B6024F029702BB0297022B0207016E00ADFFBCFEA3FE37FDF8FDD4FDD4FDD4;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h01920016FE6DFD20FCD8FDB0FF0F0080014A015C01B601EC020701EC01B60192;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hF4C3F4C3F5E3F7B7FA3FFD8C003501EC02DF036F03B703B703DB03DB03DB0303;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h07280848098C0A1C0AAC0A1C08FC0800057802970065FE13FC24F9F7F7B7F5E3;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h0138022B027301DA0031FE25FC48FA3FF8D7F88FF8D7FA87FD44002302DF0578;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFF52FFD300F00180019201C80126003AFF64FE13FCFCFC90FCB4FD68FE7FFFCA;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h057803DB02070065FF21FDD4FCD8FC24FB16FACFFB5EFC00FC48FCD8FD8CFEA3;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFDD4FCD8FC6CFCD8FDD4FF21011402DF04E9077008FC0A1C0A1C098C080006E0;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h04A103FF01A4FED9FCD8FB16F9AFF8D7F88FF88FF9AFFB16FCB4FE6DFED9FE6D;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h02730303036F0393034B03270297019200DE006500650126022B032704230459;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hFB16FCB4FEC7FFE5008000C8010201380180020701DA0180016E0180018001A4;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFF64FF7FFF76FF21FF21FED9FE5BFE13FE37FF0FFF49FE7FFCB4FA3FF9AFFA87;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h08480800065003DB0065FD20F9F7F847F847F8D7F9F7FBA6FD68FEEB00350011;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hF7B7F91FFBA6FE910114034B04A106500890098C098C08FC07B80698072807B8;
defparam sdpb_inst_0.INIT_RAM_11 = 256'hFA3FFC24FE5B00BF027303B704A10423024FFFDCFDD4FC00FA3FF91FF7B7F76F;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h0CEB0B3C08FC069805C003DB01A40053FE91FD8CFCB4FB5EF9AFF967F91FF8D7;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h034B024FFFA3FC90F91FF5E3F433F4C3F703FBA6009B04E908FC0B3C0C5B0D7B;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFDD4FDF8FDF8FD20FC6CFBA6FACFFB16FC48FC6CFCD8FDD4FEA3FFE0015C0297;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h0126FE7FFC00FA87FACFFBDCFD20FEA3FF40FF0FFEB5FF0FFF9AFF9AFEFDFE49;
defparam sdpb_inst_0.INIT_RAM_16 = 256'hF9F7FA87FC00FE5B0065024F04E908900BCC0E9B0F2B0E0B0BCC0A1C072803DB;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h011401140065FE5BFB5EF8D7F7B7F88FFBA6FEFD01B6022B00B6FEC7FCFCFB16;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h0D7B0B3C084804A10114FDD4FACFF7FFF673F673F8D7FC00FE49FFE90126014A;
defparam sdpb_inst_0.INIT_RAM_19 = 256'hF284EFB4EE94F164F553FACF002804E908900A1C0B3C0B3C0C5B0E0B0E9B0E0B;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hFFB50023006E0180032703FF053006080530036F0065FD44FBA6FA3FF88FF5E3;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h07B804A10080FB16F5E3F1F4F044F044F284F4C3F7FFFB5EFD20FE37FF91FFE5;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h02070327053008480BCC0F2B0FBB0D7B0B3C0A1C0AAC0BCC0BCC0B3C0AAC098C;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFB5EF9AFF967FA3FFB16FBA6FBA6FACFF967F7FFF673F4C3F4C3F703FACFFF0F;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h05C00207001AFF52FF6D005301A401DA0053FD8CFC24FD20FFB5027301C8FE91;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hF967F8D7F7B7F76FF7B7F88FFBA6003104E9098C0CEB0F2B104B0F2B0CEB0A1C;

endmodule //ram1_512
