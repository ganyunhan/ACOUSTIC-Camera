//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Sun Oct 09 16:33:37 2022

module ram0_512 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [8:0] ada;
input [15:0] din;
input [8:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[8:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({gw_gnd,adb[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h0073FFFBFFC4FFE9FF9A0020007C0008FFD9FF5CFFC5014A00A9FF2BFF8DFFEB;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFEFA001CFFE6FEEA0065004EFF8100CA0076FFC700F5007DFF960034FFEFFFD2;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFFE8FE97FFC400A6FF970075FF9FFE9F009C0106FFF300C500CBFF8F00AB0077;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h00C60009FF090025006CFF8F000BFFBA00B401AF00BEFEF9FF81FF3EFF26010B;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hFFB5FF5EFF5E000EFF45FEF100E10021FEE600370023FFAA007C001B00610104;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h00A6FF8CFFEF00CF004AFFC4FF26FEFB001A00F60062FF5FFFD4011B007CFFDD;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hFFF8008EFFD5FFD300A7FFDFFF270008FF7BFEFBFFD2FF21FFB200CDFF57FFB5;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFEE4FF25FEDBFF5700DAFFC8FFE9FFDCFFD50074FFBFFFE3FF50FF68007DFFEE;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h00950005FFEA00E3005DFF0EFFF2FF4EFEE0008CFF83FFD100B0FF60FFFA0035;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFFA500E3FF2CFF3500F4FF75FF6D0116FF74FF3A00AEFF3AFF09FFFEFF78FFDA;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFF10001900ABFF71FFA3FFFDFF45006A00FDFF4CFFA50094FFAFFFD9006DFF4A;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h000DFF9AFFF0006CFFF7FFDDFFBBFFA700D70076FF0600280136001F00320018;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFFD0FFF5FFAB001F002C001600C400C300810058FFC8FF72FFCFFFB7FF9A0018;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h00460039FFC3002C002CFFD90069005C0002005C0032FFF7003D003CFF92FF44;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h00160038FFB8FF61006F00A0FFC1FFDC0049004500810027FF56FFEC00720001;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h001AFF6BFF55FFD80013009A00F20008FFA40049003800730061FF27FF7D003A;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h00130062001A0001000100D30139002EFFC8007500880016FFABFF47FF41FFE2;
defparam sdpb_inst_0.INIT_RAM_11 = 256'hFFBD001F002C005900BD005800A10141006DFFD40009FFFA007C0074FEFAFEC4;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFE6FFF4004EFFDEFF980069006DFFB1FFFA00D700E40052FF9AFF7F00390023;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hFFE9FF68FF4CFFB70031FFEAFFACFFDF004000BB006FFFCC005D00DF0054FFFE;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h001BFFADFEF0FF41FF3DFF4700380026FF9A005300BA008E009E0026000D0059;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h00190004FF62FEF6FFECFFCAFF35FFA0FFB20016012800FD0071009B0038FFD1;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h00D80058FF09FF4F003C00E400E9FF87FF17004100AF0095000FFF42FFF2009C;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hFFB6FFA400AE00C70042000EFF78FF80FFCCFF78002400A1FFAFFF91FFF1001F;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h00050056003BFF17FF5D00A900B3005BFFE6FFC00053FFF4FF3AFFBA008A0084;
defparam sdpb_inst_0.INIT_RAM_19 = 256'hFF4BFF0E00270082002FFF89FF22002600DFFFF5FF46FFCB007B0036FF9EFFC9;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h0036FF3FFFC20042FFE00011000FFFB3FFFD0040FFE2FFEA003D00160060007F;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hFFC5007100290019003EFFB4FFB6FFF0FFC00064006BFF50FFA7002DFFBC0047;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h0051FF78FF76003200380017FFEE001A009E0004FF6DFFE90001FFF00006FF96;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFF61FFC4FFF200020092002CFFC4007F003AFF7C00090028FFB9FFD8FFD50027;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h0008FFAF00C6003AFF5700930055FF930079FFC1FF3700A1FFF4FEBAFFB9FFFB;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h00D100B9004A0041000FFFBCFFB3FFC5FFD7FFE0FF7EFF2DFFD90003FF970032;

endmodule //ram0_512
