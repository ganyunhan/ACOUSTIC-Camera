//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Tue Sep 27 23:11:56 2022

module ram0_512 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [8:0] ada;
input [15:0] din;
input [8:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[8:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({gw_gnd,adb[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFF22FF1EFF45FF7AFF8DFFADFFCEFFE000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h029B027F02360227023001FC01BB01B6019D0168010D008600660040FFC1FF45;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFF8DFF45FEA4FE35FE4DFE28FE2CFDB7FCF2FCC6FD62FE44FFC00173027802C1;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h00D2FFF7FED0FE42FE06FDD6FDD5FDD4FDBDFD8CFDA8FDE0FE8BFF3FFFB9FFD4;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h0139015601A201E6020301F701BF019801A20231029002B302AB023A02120197;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h02BC035303B403B203D703D903E4034301DD0066FEC2FD52FCCEFD73FEC5003A;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h0619031600D8FE85FC85FA70F823F637F4E8F4ABF596F74FF9A7FCE3FFC401A3;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hF904F891F8B5FA0EFCB2FF90025604FB06EC0804095A0A010A990A56092A0848;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFF9BFE58FD28FC98FCA4FD37FE45FF8000F502070274020E0098FE89FCABFAA6;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFB49FAC4FB3BFBE7FC3AFCB5FD64FE67FF41FFA800B90175018B01C5015B0060;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h0464070408B209F90A2709BF0851071305CD042D026A00ACFF63FE15FCFFFC50;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hF899F87EF961FAD4FC52FE29FEDEFE87FDFAFD0BFC6BFCB7FD98FED600A40290;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h00FD0076005700F101FC02ED04000452049504450236FF5BFD34FB6EF9ECF8F4;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h016901F301F20189017001790186018B024802ED035A03970359032D02C501C2;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFE1FFEE2FF58FEB6FD2DFAA9F999FA60FAF1FC45FE6EFFBA006800BD00F50130;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hF839F8AEF9B2FB46FD17FE9B00090035FF79FF71FF86FF2BFF21FEF1FE71FE1D;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h08310972099B0922080A06AE06FC07A2082B083406B50472011BFDC4FA8EF86E;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h02BF005BFE2DFC68FA85F960F7F2F768F79EF8B6FB18FDFD009C02E3046B05DC;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFEE4FDB3FCE6FBB4F9F3F95EF942F8C3F9E1FBC1FDDF004D022B03770487045E;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hF660FA96FFB2040908440AF20C1D0D560D300B97098506F305E7046101F700A0;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFC19FC72FCACFDA7FE75FF960112025F033D02B0003AFD36F9D3F678F458F485;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hFF39FF21FEBFFEEDFF89FFA7FF26FE68FDE4FDE5FE0FFD4EFC8DFBD4FAF0FAE4;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h0B240E300F380E660C3A0A7807E1047001B2FF04FC79FAACFAA6FBA3FCD6FE5E;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hFAEFFE5C0145024F010DFF30FD51FB7FFA04FA5BFB98FDE6FFFF01ED043F07DB;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hF6A4F649F832FB6EFDE4FF9D00F601590115011C009FFEE2FBFAF941F7CFF830;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h081309D10B200B340C070DBE0EA40E220DB20BCA08EA056601C0FE77FB68F87F;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h057303DE0119FDC7FBE7FA8FF8EEF68BF327F03AEE7DF0A2F47AF996FF3503ED;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hF200F44EF73CFAD1FCE0FDF9FF53FFF1FFAF000D005B012E02E003D904E60601;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h0BA20A300A770B9C0BE90B4F0AD809CA0836054E0177FC31F6E3F28CF07CF010;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hF9BBF83CF6D6F500F499F661F9FEFE3601A602EB04AB079D0B100E9B0FF10DFD;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h00CDFE13FC3AFCC5FF180211023DFF41FBF0F9DFF961FA02FAFAFB88FBC0FB01;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h0405089D0C6C0EB710480F820D6D0AC206B80294006CFF5DFF61000B017201EB;

endmodule //ram0_512
