//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.08
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Sat Oct 22 12:44:23 2022

module ram2_512 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [8:0] ada;
input [15:0] din;
input [8:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[8:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({gw_gnd,adb[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFF7FFF2CFF1FFF28FF63FF84FF99FFBFFFD7FFEC000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h02B202B00292025F02230230022001D801B401B20184014900C9006B0060000D;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFFD7FFB7FF6FFF08FE58FE40FE3FFE27FE0FFD54FCC2FCFCFDC4FEDA00980202;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h01EE0138007AFF6BFE76FE29FDE8FDD4FDD3FDD2FD9FFD93FDBBFE21FEE8FF7D;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hFF7100CF0153016C01CC01F3020801DC01AC018E01D9026E029E02C002770220;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h00BA023F0306038E03B503C103DC03E003BE02A60132FFAAFE04FCF0FCF8FE06;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h08C7078404A501FFFFC9FD89FBA0F959F732F581F4A6F4F5F651F848FB13FE5B;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFBC3F9C3F8B0F891F91CFB33FE0400E00391060B076D08A709BD0A440AAE09C8;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h00DF000CFF13FDBEFCCEFC8FFCD3FDAEFECD002D0187025002630184FFA5FDA8;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFCACFBE2FAE5FAE9FB8EFC19FC63FD06FDCAFEE8FF650018012C018601A201BB;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h01A0034905A107E7095B0A320A09093307A40695050A036A018B000EFECAFD85;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hF967F8BBF882F8BBFA15FB71FD38FEADFEC6FE4BFD99FCA1FC7AFD0CFE25FF8F;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h0252015B00B800560084016F02660375043E046704A0038600E0FE41FC61FAAB;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h0113014301A5021201B90179016D0188017901D202A3031F03850385033D0316;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFE43FE0CFE65FF3DFF27FE28FC08F9D8F9E2FAADFB5CFD4CFF280015009900D5;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hF94DF82FF860F915FA59FC25FDCDFF530054FFDBFF5AFF8DFF5CFF1CFF1BFEB6;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h04EF06F408F309A0097008BF074D069E075B07D8085F07A505C50302FF80FC48;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h04AA03C101B2FF3FFD63FB79F9F3F8BEF783F77BF7EDF9B7FC66FF4801AF03BF;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h014CFFE0FE36FD5AFC6DFAE5F974F96EF8EEF911FABCFCABFF00014502CA0406;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hF42AF52AF803FD0901BC060D09C90B8A0CB20D8C0C820ABE0843064605750329;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFAB7FB6AFC6DFC6DFD1CFE09FEE8004401B702DA034101B5FEDDFBB1F837F53B;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hFD87FEEBFF3FFEF4FEB6FF3DFFA8FF80FEC8FE24FDCBFE0FFDCAFCEBFC3FFB69;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h05DA096E0CA50EFB0F050D7D0B500988063603230071FDD3FB74FA74FB0EFC29;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hF7B5F933FC93FFC9022001DF003EFE43FC8AFA9BFA04FACAFC9AFEEA00E802D7;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hFA07F770F648F6D6F9B7FCAEFEC2004801500132011900FE0003FD9CFA9DF864;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h015C061F090B0A800B450B600CD10E5D0E7A0DF50D110A7D076603A50037FD05;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h058C05F304D002C6FF79FCB8FB52F9D4F802F4FDF1BCEF1AEEFDF264F68FFC5C;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hF00FF0B4F324F572F8FEFBF9FD69FE90FFCEFFCCFFCB003A009501F60370043A;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h0F460CD70AC80A1E0AFA0BF30B9E0B250A67093206FF03B2FF25F9AEF4A8F156;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFB78FA83F8FBF7ADF5EEF492F51FF7EDFBE500130262038A05EE092B0CC10FB5;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h01D101A8FF9EFCF6FC30FDAE008902B30109FDADFABCF984F983FA8AFB38FBC4;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hFCAB018206140AA90D810FB110290EA90C400923048E016DFFC2FF51FF8A00B8;

endmodule //ram2_512
