//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Wed Sep 28 20:31:39 2022

module acos_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [23:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h787B7D808285878A8C8F9295989B9EA1A4A7ABAFB2B6BBBFC4C9CED4DBE3EE08;
defparam prom_inst_0.INIT_RAM_01 = 256'h3B3D3E4042434547494A4C4E5052535557595B5D5F61636567696B6D6F727476;
defparam prom_inst_0.INIT_RAM_02 = 256'h0C0D0E10111214151718191B1C1E1F2122242527282A2B2D2E30313335363839;
defparam prom_inst_0.INIT_RAM_03 = 256'hE4E5E6E7E8E9EBECEDEEEFF1F2F3F4F6F7F8F9FBFCFDFF00010204050608090A;
defparam prom_inst_0.INIT_RAM_04 = 256'hC0C1C2C3C4C5C6C7C8CACBCCCDCECFD0D1D2D3D5D6D7D8D9DADBDDDEDFE0E1E2;
defparam prom_inst_0.INIT_RAM_05 = 256'h9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B9BABBBCBDBEBF;
defparam prom_inst_0.INIT_RAM_06 = 256'h8182838485868788898A8A8B8C8D8E8F909192939495969798999A9B9C9C9D9E;
defparam prom_inst_0.INIT_RAM_07 = 256'h6566676868696A6B6C6D6E6F6F70717273747576767778797A7B7C7D7E7F7F80;
defparam prom_inst_0.INIT_RAM_08 = 256'h4A4B4C4D4D4E4F5051525253545556575758595A5B5C5C5D5E5F606162626364;
defparam prom_inst_0.INIT_RAM_09 = 256'h3131323334353536373838393A3B3C3C3D3E3F40404142434444454647484949;
defparam prom_inst_0.INIT_RAM_0A = 256'h18191A1A1B1C1D1D1E1F202021222323242526272728292A2A2B2C2D2D2E2F30;
defparam prom_inst_0.INIT_RAM_0B = 256'h000102030304050506070808090A0B0B0C0D0E0E0F1011111213141415161717;
defparam prom_inst_0.INIT_RAM_0C = 256'hE9EAEBECECEDEEEEEFF0F0F1F2F3F3F4F5F5F6F7F8F8F9FAFBFBFCFDFDFEFF00;
defparam prom_inst_0.INIT_RAM_0D = 256'hD3D4D4D5D6D7D7D8D9D9DADBDBDCDDDDDEDFE0E0E1E2E2E3E4E4E5E6E7E7E8E9;
defparam prom_inst_0.INIT_RAM_0E = 256'hBDBEBFBFC0C1C1C2C3C3C4C5C5C6C7C7C8C9C9CACBCCCCCDCECECFD0D0D1D2D2;
defparam prom_inst_0.INIT_RAM_0F = 256'hA8A9A9AAABABACADADAEAFAFB0B1B1B2B3B3B4B5B5B6B7B7B8B9B9BABBBBBCBD;
defparam prom_inst_0.INIT_RAM_10 = 256'h939495959696979898999A9A9B9C9C9D9E9E9FA0A0A1A2A2A3A3A4A5A5A6A7A7;
defparam prom_inst_0.INIT_RAM_11 = 256'h7F7F8081818283838485858686878888898A8A8B8C8C8D8D8E8F8F9091919293;
defparam prom_inst_0.INIT_RAM_12 = 256'h6B6B6C6D6D6E6E6F707071727273737475757677777879797A7A7B7C7C7D7E7E;
defparam prom_inst_0.INIT_RAM_13 = 256'h57585859595A5B5B5C5C5D5E5E5F60606161626363646565666667686869696A;
defparam prom_inst_0.INIT_RAM_14 = 256'h43444545464647484849494A4B4B4C4D4D4E4E4F505051515253535454555656;
defparam prom_inst_0.INIT_RAM_15 = 256'h303131323233343435353637373838393A3A3B3C3C3D3D3E3F3F404041424243;
defparam prom_inst_0.INIT_RAM_16 = 256'h1D1E1E1F1F20212122222324242525262627282829292A2B2B2C2C2D2E2E2F2F;
defparam prom_inst_0.INIT_RAM_17 = 256'h0A0B0B0C0C0D0E0E0F0F10111112121313141515161617181819191A1B1B1C1C;
defparam prom_inst_0.INIT_RAM_18 = 256'hF7F8F8F9FAFAFBFBFCFCFDFEFEFFFF0001010202030404050506060708080909;
defparam prom_inst_0.INIT_RAM_19 = 256'hE5E5E6E6E7E7E8E9E9EAEAEBECECEDEDEEEEEFF0F0F1F1F2F3F3F4F4F5F5F6F7;
defparam prom_inst_0.INIT_RAM_1A = 256'hD2D3D3D4D4D5D5D6D7D7D8D8D9DADADBDBDCDCDDDEDEDFDFE0E0E1E2E2E3E3E4;
defparam prom_inst_0.INIT_RAM_1B = 256'hC0C0C1C1C2C2C3C4C4C5C5C6C6C7C8C8C9C9CACACBCCCCCDCDCECFCFD0D0D1D1;
defparam prom_inst_0.INIT_RAM_1C = 256'hADAEAEAFAFB0B1B1B2B2B3B3B4B5B5B6B6B7B7B8B9B9BABABBBBBCBDBDBEBEBF;
defparam prom_inst_0.INIT_RAM_1D = 256'h9B9B9C9C9D9E9E9F9FA0A0A1A2A2A3A3A4A4A5A6A6A7A7A8A8A9AAAAABABACAD;
defparam prom_inst_0.INIT_RAM_1E = 256'h88898A8A8B8B8C8C8D8E8E8F8F90909192929393949495969697979898999A9A;
defparam prom_inst_0.INIT_RAM_1F = 256'h767777787879797A7B7B7C7C7D7D7E7F7F808081818283838484858686878788;
defparam prom_inst_0.INIT_RAM_20 = 256'h64646565666767686869696A6B6B6C6C6D6D6E6F6F7070717172737374747575;
defparam prom_inst_0.INIT_RAM_21 = 256'h5152525354545555565657585859595A5A5B5C5C5D5D5E5F5F60606161626363;
defparam prom_inst_0.INIT_RAM_22 = 256'h3F3F40414142424343444545464647474849494A4A4B4C4C4D4D4E4E4F505051;
defparam prom_inst_0.INIT_RAM_23 = 256'h2C2D2D2E2F2F30303132323333343435363637373838393A3A3B3B3C3D3D3E3E;
defparam prom_inst_0.INIT_RAM_24 = 256'h1A1A1B1B1C1D1D1E1E1F2020212122222324242525262727282829292A2B2B2C;
defparam prom_inst_0.INIT_RAM_25 = 256'h07080809090A0B0B0C0C0D0D0E0F0F1010111212131314141516161717181919;
defparam prom_inst_0.INIT_RAM_26 = 256'hF4F5F5F6F6F7F8F8F9F9FAFBFBFCFCFDFEFEFFFF000101020203030405050606;
defparam prom_inst_0.INIT_RAM_27 = 256'hE1E2E2E3E3E4E5E5E6E6E7E8E8E9E9EAEBEBECECEDEEEEEFEFF0F1F1F2F2F3F4;
defparam prom_inst_0.INIT_RAM_28 = 256'hCECFCFD0D0D1D2D2D3D3D4D5D5D6D6D7D8D8D9D9DADBDBDCDCDDDEDEDFDFE0E1;
defparam prom_inst_0.INIT_RAM_29 = 256'hBABBBCBCBDBEBEBFBFC0C1C1C2C2C3C4C4C5C5C6C7C7C8C8C9CACACBCBCCCDCD;
defparam prom_inst_0.INIT_RAM_2A = 256'hA7A7A8A9A9AAABABACACADAEAEAFAFB0B1B1B2B3B3B4B4B5B6B6B7B7B8B9B9BA;
defparam prom_inst_0.INIT_RAM_2B = 256'h93949495959697979899999A9A9B9C9C9D9E9E9F9FA0A1A1A2A2A3A4A4A5A6A6;
defparam prom_inst_0.INIT_RAM_2C = 256'h7F7F808181828283848485868687888889898A8B8B8C8D8D8E8E8F9090919292;
defparam prom_inst_0.INIT_RAM_2D = 256'h6A6B6B6C6D6D6E6F6F7071717272737474757676777878797A7A7B7B7C7D7D7E;
defparam prom_inst_0.INIT_RAM_2E = 256'h555656575858595A5A5B5C5C5D5E5E5F60606162626364646565666767686969;
defparam prom_inst_0.INIT_RAM_2F = 256'h4040414242434444454646474848494A4A4B4C4C4D4E4E4F5050515252535454;
defparam prom_inst_0.INIT_RAM_30 = 256'h2A2A2B2C2C2D2E2E2F3030313233333435353637373839393A3B3B3C3D3E3E3F;
defparam prom_inst_0.INIT_RAM_31 = 256'h131414151617171819191A1B1B1C1D1E1E1F2020212223232425252627272829;
defparam prom_inst_0.INIT_RAM_32 = 256'hFCFCFDFEFFFF000102020304040506070708090A0A0B0C0C0D0E0F0F10111212;
defparam prom_inst_0.INIT_RAM_33 = 256'hE4E4E5E6E7E7E8E9EAEAEBECEDEDEEEFF0F0F1F2F3F3F4F5F6F6F7F8F9F9FAFB;
defparam prom_inst_0.INIT_RAM_34 = 256'hCBCBCCCDCECFCFD0D1D2D2D3D4D5D6D6D7D8D9DADADBDCDDDDDEDFE0E0E1E2E3;
defparam prom_inst_0.INIT_RAM_35 = 256'hB0B1B2B3B4B5B5B6B7B8B9BABABBBCBDBEBEBFC0C1C2C3C3C4C5C6C7C7C8C9CA;
defparam prom_inst_0.INIT_RAM_36 = 256'h9596979898999A9B9C9D9E9F9FA0A1A2A3A4A5A5A6A7A8A9AAABABACADAEAFB0;
defparam prom_inst_0.INIT_RAM_37 = 256'h78797A7B7C7D7D7E7F80818283848586878888898A8B8C8D8E8F909191929394;
defparam prom_inst_0.INIT_RAM_38 = 256'h595A5B5C5D5E5F606162636465666768696A6B6B6C6D6E6F7071727374757677;
defparam prom_inst_0.INIT_RAM_39 = 256'h3738393A3B3C3D3F404142434445464748494A4B4C4D4E505152535455565758;
defparam prom_inst_0.INIT_RAM_3A = 256'h111314151618191A1B1C1E1F2021222325262728292A2C2D2E2F303132343536;
defparam prom_inst_0.INIT_RAM_3B = 256'hE6E8E9EBECEEEFF0F2F3F5F6F7F9FAFBFDFEFF010203050607080A0B0C0E0F10;
defparam prom_inst_0.INIT_RAM_3C = 256'hB2B4B5B7B9BBBDBEC0C2C4C5C7C9CACCCECFD1D2D4D6D7D9DADCDDDFE0E2E3E5;
defparam prom_inst_0.INIT_RAM_3D = 256'h66696C6F7275787B7D808285878A8C8F919395989A9C9EA0A2A4A6A8AAACAEB0;
defparam prom_inst_0.INIT_RAM_3E = 256'h000000000000000000000000000000000019242C33393E43484C5155585C6063;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0606060606060606060606060606060606060606060606060606060606060607;
defparam prom_inst_1.INIT_RAM_01 = 256'h0606060606060606060606060606060606060606060606060606060606060606;
defparam prom_inst_1.INIT_RAM_02 = 256'h0606060606060606060606060606060606060606060606060606060606060606;
defparam prom_inst_1.INIT_RAM_03 = 256'h0505050505050505050505050505050505050505050505060606060606060606;
defparam prom_inst_1.INIT_RAM_04 = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam prom_inst_1.INIT_RAM_05 = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam prom_inst_1.INIT_RAM_06 = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam prom_inst_1.INIT_RAM_07 = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam prom_inst_1.INIT_RAM_08 = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam prom_inst_1.INIT_RAM_09 = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam prom_inst_1.INIT_RAM_0A = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam prom_inst_1.INIT_RAM_0B = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam prom_inst_1.INIT_RAM_0C = 256'h0404040404040404040404040404040404040404040404040404040404040405;
defparam prom_inst_1.INIT_RAM_0D = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_0E = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_0F = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_10 = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_11 = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_12 = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_13 = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_14 = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_15 = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_16 = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_17 = 256'h0404040404040404040404040404040404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_18 = 256'h0303030303030303030303030303030404040404040404040404040404040404;
defparam prom_inst_1.INIT_RAM_19 = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_1A = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_1B = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_1C = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_1D = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_1E = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_1F = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_20 = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_21 = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_22 = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_23 = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_24 = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_25 = 256'h0303030303030303030303030303030303030303030303030303030303030303;
defparam prom_inst_1.INIT_RAM_26 = 256'h0202020202020202020202020202020202020202030303030303030303030303;
defparam prom_inst_1.INIT_RAM_27 = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_28 = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_29 = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_2A = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_2B = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_2C = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_2D = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_2E = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_2F = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_30 = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_31 = 256'h0202020202020202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_32 = 256'h0101010101010202020202020202020202020202020202020202020202020202;
defparam prom_inst_1.INIT_RAM_33 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam prom_inst_1.INIT_RAM_34 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam prom_inst_1.INIT_RAM_35 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam prom_inst_1.INIT_RAM_36 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam prom_inst_1.INIT_RAM_37 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam prom_inst_1.INIT_RAM_38 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam prom_inst_1.INIT_RAM_39 = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam prom_inst_1.INIT_RAM_3A = 256'h0101010101010101010101010101010101010101010101010101010101010101;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000001010101010101010101010101;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //acos_rom
