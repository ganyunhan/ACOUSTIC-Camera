//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.08
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Created Time: Thu Oct 13 17:53:14 2022

module ram0_512 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [8:0] ada;
input [15:0] din;
input [8:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[8:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({gw_gnd,adb[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFFC5FFE2FFFFFFFCFFF4FFF3FFF3FFF2FFE2FFCAFFBEFFE2FFE8000F00490018;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFFFBFFCE0005003B00040015000AFFBAFFB2FFB7FFC800180013FFF900260008;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h001C000DFFF10005FFE2FFFAFFFC0023FFDCFFAE0006FF68FF89FFFBFFA5FFD6;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hFFBEFFC9FFE9FFA3FFFC0053000AFFE6002AFFEEFFA30000000800120068003B;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h004DFFFF000BFFFFFFBBFFCAFFBDFF7CFFB0FFEFFFC0FFD80033FFF7FFE4002F;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hFFFE00050005FFF6FFE500090019FFEAFFD7FFF20002FFE9FFE70002FFE0001B;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hFFC4FFCEFFF50019002E0025FFFFFFD6FFD5FFDFFFE6FFF6FFE6FFFCFFF9FFF2;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h001800230021FFDBFFCCFFD9FFC7FFFA001D000F002E0014FFF50020FFFFFFC9;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFFAEFFC9FFEF00290016FFFE00380021FFDFFFCEFF96FF9EFFE6FFEE00040032;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFFE8FFEAFFEDFFD9FFDDFFD8FFFB002A001CFFFE0000000C00150018FFEBFFAA;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h00040002FFA3FFD9FFF4FFB700020010FFF800270024FFF8FFF7FFE2FFE8FFFA;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hFFEB000A004B0022000E000BFFCBFFE90013FFC8FFD80013000000240035FFE6;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFFF4FFD6FFDDFFF7FFFF0018001D0011000C0000FFD7FFBEFFF4FFE4FFD6FFF7;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hFFD4FFF8FFECFFD00015FFFAFFD9000DFFE0FFCD0001FFDCFFEF00290004FFEB;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h0003FFFCFFEFFFFF0001FFF80017FFF7FFE20008000400100029FFF500010009;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hFFE9FFCEFFDDFFD4FFC6FFF1FFF7FFDBFFFF000200060018FFF1FFEE0025000E;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h0017FFF7FFD7FFF6FFECFFDDFFDEFFCFFFCE0000002400240039002BFFF3FFEC;
defparam sdpb_inst_0.INIT_RAM_11 = 256'hFFE2FFFCFFFAFFEEFFFCFFDCFFD800130019FFF3FFF6FFF7FFE800180021FFFF;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFECFFE0FFEAFFF2FFFB0001FFEDFFFB00020003001E002E001A000B00150002;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h0002FFF5001B00190017001BFFF9000C002B002C0019FFFDFFF90014FFF6FFE8;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFFF90020000FFFF4001D0008FFDE000E000D00240042000200060010FFD5FFEA;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h0038005900390010001A000E000E0013FFEBFFFC00140007000600190028000E;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h0034001C002B0003FFF3001B001500010002FFF0FFFF0015FFF8FFE50000001B;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h002E001A00060023FFDFFFCCFFF9FFE4FFFE0015FFEC0012004600270023004C;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h00170022FFF4FFFCFFE0FFD90006FFFF0000000C000C001E002200240000FFF1;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h001400030004FFFFFFE8FFECFFD5FFE20000FFE2FFFA001FFFF2FFFDFFF8FFD8;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hFFF3FFD5FFC0FFF400010002000FFFFFFFEEFFEBFFF30009000D0003FFF8000B;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h00160014FFF800060017FFF3FFF30001FFF7000DFFFCFFF0002200350013FFF7;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hFFFE00240006FFE900130010FFF9FFD7FFC4FFF000200000FFECFFFC00080003;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFFE5000B000100050001FFD3FFFD0016001B002F001D00180006FFD7FFF3FFFC;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h00390025FFF6001C00230008001E001000200026FFECFFDEFFDFFFCCFFFBFFF7;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h000700010001FFE2FFF00009FFFA0007FFFEFFD4FFECFFEDFFDE001200210011;

endmodule //ram0_512
